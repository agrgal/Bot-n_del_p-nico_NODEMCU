NodeMCU_EMISOR_V01

.TRAN 1ms 100ms
* .AC DEC 100 100 1MEG
.END
